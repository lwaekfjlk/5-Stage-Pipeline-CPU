`timescale 1ns / 1ps

`define DEBUG

`ifdef XILINX_ISIM
	`define SIMULATING
`endif
